`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/11/2024 09:25:38 PM
// Design Name: 
// Module Name: quadSevenSeg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module quadSevenSeg(
    output [6:0] seg,
    output dp,
    output an0,
    output an1,
    output an2,
    output an3,
    input [7:0] char0, 
    input [7:0] char1,
    input [7:0] char2,
    input [7:0] char3, 
    input clk
    );
    
    reg [7:0] hexIn;
    reg [1:0] ns; // next stage
    reg [1:0] ps; // present stage
    reg [3:0] dispEn; // which 7seg is active
    wire [6:0] segments;
    assign seg=segments;
    hexTo7Segment segDecode(segments,hexIn);
    assign dp=1;
    assign {an3,an2,an1,an0}=~dispEn;


    always @(posedge clk)
        ps=ns;

    always @(ps) 
        ns=ps+1;
    
    always @(ps)
        case(ps)
            2'b00: dispEn=4'b0001;
            2'b01: dispEn=4'b0010;
            2'b10: dispEn=4'b0100;
            2'b11: dispEn=4'b1000;
        endcase
    
    always @(ps)
        case(ps)
            2'b00: hexIn=char0;
            2'b01: hexIn=char1;
            2'b10: hexIn=char2;
            2'b11: hexIn=char3;
        endcase

    
endmodule
